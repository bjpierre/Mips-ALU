---- 5 to 32 dec---
library IEEE;
use IEEE.std_logic_1164.all;
entity bitdecoder is
	port(bitin : in std_logic_vector(4 downto 0);
	     bitout : out std_logic_vector(31 downto 0);
	     wen : in std_logic);
end bitdecoder;

architecture Behavioral of bitdecoder is

begin
process(bitin,wen)
begin
	
	if(wen = '0') then
		bitout <= "00000000000000000000000000000000";
	else
		case bitin is 
			when "00000" => bitout <= "00000000000000000000000000000001";
			when "00001" => bitout <= "00000000000000000000000000000010";
			when "00010" => bitout <= "00000000000000000000000000000100";
			when "00011" => bitout <= "00000000000000000000000000001000";
			when "00100" => bitout <= "00000000000000000000000000010000";
			when "00101" => bitout <= "00000000000000000000000000100000";
			when "00110" => bitout <= "00000000000000000000000001000000";
			when "00111" => bitout <= "00000000000000000000000010000000";
			when "01000" => bitout <= "00000000000000000000000100000000";
			when "01001" => bitout <= "00000000000000000000001000000000";
			when "01010" => bitout <= "00000000000000000000010000000000";
			when "01011" => bitout <= "00000000000000000000100000000000";
			when "01100" => bitout <= "00000000000000000001000000000000";
			when "01101" => bitout <= "00000000000000000010000000000000";
			when "01110" => bitout <= "00000000000000000100000000000000";
			when "01111" => bitout <= "00000000000000001000000000000000";
			when "10000" => bitout <= "00000000000000010000000000000000";
			when "10001" => bitout <= "00000000000000100000000000000000";
			when "10010" => bitout <= "00000000000001000000000000000000";
			when "10011" => bitout <= "00000000000010000000000000000000";
			when "10100" => bitout <= "00000000000100000000000000000000";
			when "10101" => bitout <= "00000000001000000000000000000000";
			when "10110" => bitout <= "00000000010000000000000000000000";
			when "10111" => bitout <= "00000000100000000000000000000000";
			when "11000" => bitout <= "00000001000000000000000000000000";
			when "11001" => bitout <= "00000010000000000000000000000000";
			when "11010" => bitout <= "00000100000000000000000000000000";
			when "11011" => bitout <= "00001000000000000000000000000000";
			when "11100" => bitout <= "00010000000000000000000000000000";
			when "11101" => bitout <= "00100000000000000000000000000000";
			when "11110" => bitout <= "01000000000000000000000000000000";
			when "11111" => bitout <= "10000000000000000000000000000000";
			when others => bitout <= "00000000000000000000000000000000";
		end case;
	end if;
end process;
end Behavioral;
